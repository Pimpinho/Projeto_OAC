// COMPILE: iverilog.exe -g2012 -o riscvsingle_p1.vcd -tvvp .\riscvsingle_p1.sv
// SIMULATE: vvp riscvsingle_p1
// https://www.edaplayground.com/

module testbench();

  logic        clk;
  logic        reset;

  logic [31:0] WriteData, DataAdr;
  logic        MemWrite;

  // instantiate device to be tested
  top dut(clk, reset, WriteData, DataAdr, MemWrite, PCSrc);
  
  // initialize test
  initial
    begin
      reset <= 1; # 22; reset <= 0;
    end

  // generate clock to sequence tests
  always
    begin
      clk <= 1; # 5; clk <= 0; # 5;
    end

  // check results
  always @(negedge clk)
    begin
      if(MemWrite) begin
        if(DataAdr === 100 & WriteData === 25) begin
          $display("Simulation succeeded");
          $stop;
        end else if (DataAdr !== 96) begin
          $display("Simulation failed");
          $stop;
        end
      end
    end
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module top(input  logic        clk, reset, 
           output logic [31:0] WriteData, DataAdr, 
           output logic        MemWrite,
           output logic        PCSrc);  //// [MODIFICAÇAO] PCSrc nao estava sendo passado como saida do modulo e era exigido no testbench
                                        //// como esta na saida do moulo mais acima, agora esta visivel para os outros niveis ////

  logic [31:0] PC, Instr, ReadData;
  
  // instantiate processor and memories
  riscvsingle rvsingle(clk, reset, PC, Instr, MemWrite, DataAdr, 
                     WriteData, ReadData, PCSrc); //// [MODIFICAÇAO] PCSrc nao estava sendo passado ////
                                                  
  imem imem(PC, Instr);
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module riscvsingle(input  logic        clk, reset,
                  output logic [31:0] PC,
                  input  logic [31:0] Instr,
                  output logic        MemWrite,
                  output logic [31:0] ALUResult, WriteData,
                  input  logic [31:0] ReadData,
                  output logic        PCSrc); //// [MODIFICAÇAO] antes o PCSrc nao estava sendo passado como saida do modulo
                                              //// logo nao se tornava visivel para outros modulos ////

  logic       ALUSrc, RegWrite, Jump, Zero;   //// [MODIFICAÇAO] PCSrc foi removido dessa declaracao e foi para a saida do modulo ////
  logic [1:0] ResultSrc, ImmSrc;
  logic [2:0] ALUControl;

  controller c(Instr[6:0], Instr[14:12], Instr[30], Zero,
               ResultSrc, MemWrite, PCSrc,
               ALUSrc, RegWrite, Jump,
               ImmSrc, ALUControl);
  datapath dp(clk, reset, ResultSrc, PCSrc,
              ALUSrc, RegWrite,
              ImmSrc, ALUControl,
              Zero, PC, Instr,
              ALUResult, WriteData, ReadData);
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module controller(input  logic [6:0] op,
                  input  logic [2:0] funct3,
                  input  logic       funct7b5,
                  input  logic       Zero,
                  output logic [1:0] ResultSrc,
                  output logic       MemWrite,
                  output logic       PCSrc, ALUSrc,
                  output logic       RegWrite, Jump,
                  output logic [1:0] ImmSrc,
                  output logic [2:0] ALUControl);

  logic [1:0] ALUOp;
  logic       Branch;

  maindec md(op, ResultSrc, MemWrite, Branch, ALUSrc, RegWrite, Jump, ImmSrc, ALUOp);
  
  aludec ad(op[5], funct3, funct7b5, ALUOp, ALUControl);

  assign PCSrc = (Branch & Zero) | Jump; //// [MODIFICAÇAO] antes o assign era PCSrc = Branch & Zero
                                         ////Ou seja, instruçoes de Jump nao eram tratadas ////
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module maindec(input  logic [6:0] op,
              output logic [1:0] ResultSrc,
              output logic       MemWrite,
              output logic       Branch,
              output logic       ALUSrc,
              output logic       RegWrite,
              output logic       Jump,
              output logic [1:0] ImmSrc,
              output logic [1:0] ALUOp);

  logic [10:0] controls;

  assign {RegWrite, ImmSrc, ALUSrc, MemWrite,
          ResultSrc, Branch, ALUOp, Jump} = controls; //// [MODIFICAÇAO]             
  

  
  always_comb
    case(op)
    // RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
      7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
      7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
      7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type 
      7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
      7'b0010011: controls = 11'b1_00_1_0_00_0_00_0; // I-type ALU (addi, ori, andi, slti) //// [MODIFICAÇAO] antes nao existia essa linha ////
      7'b1101111: controls = 11'b1_11_0_0_10_0_00_1; // jal  //// [MODIFICAÇAO] antes nao existia essa linha ////
      default:    controls = 11'bx_xx_x_x_xx_x_xx_x; // non-implemented instruction
    endcase
endmodule

  
  // [MODIFICAÇÃO] Adicionado suporte a:
  // 1. assign de Jump em controls - para instruçoes JAL
  // 2. I-type (0010011) - operaçoes imediatas
  // 3. JAL (1101111) - jump and link
  // Controles atualizados: {RegWrite,ImmSrc,ALUSrc,MemWrite,ResultSrc,Branch,ALUOp,Jump}

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module aludec(input  logic       opb5,
             input  logic [2:0] funct3,
             input  logic       funct7b5,
             input  logic [1:0] ALUOp,
             output logic [2:0] ALUControl);

  logic  RtypeSub;
  assign RtypeSub = funct7b5 & opb5;  // TRUE for R-type subtract instruction

  always_comb
    case(ALUOp)
      2'b00:                ALUControl = 3'b000; // addition
      2'b01:                ALUControl = 3'b001; // subtraction
      default: case(funct3) // R-type or I-type ALU
                 3'b000:  if (RtypeSub) 
                            ALUControl = 3'b001; // sub
                          else          
                            ALUControl = 3'b000; // add, addi
                 3'b010:    ALUControl = 3'b101; // slt, slti
                 3'b110:    ALUControl = 3'b011; // or, ori
                 3'b111:    ALUControl = 3'b010; // and, andi
                 default:   ALUControl = 3'bxxx; // ???
               endcase
    endcase
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module datapath(input  logic        clk, reset,
               input  logic [1:0]  ResultSrc,
               input  logic        PCSrc,
               input  logic        ALUSrc,
               input  logic        RegWrite,
               input  logic [1:0]  ImmSrc,
               input  logic [2:0]  ALUControl,
               output logic        Zero,
               output logic [31:0] PC,
               input  logic [31:0] Instr,
               output logic [31:0] ALUResult,
               output logic [31:0] WriteData,
               input  logic [31:0] ReadData);

  logic [31:0] PCNext, PCPlus4, PCTarget;
  logic [31:0] ImmExt;
  logic [31:0] SrcA, SrcB;
  logic [31:0] Result;

  // PC logic
  flopr #(32) pc_reg(clk, reset, PCNext, PC);
  adder       pcadd4(PC, 32'd4, PCPlus4);
  adder       pcaddbranch(PC, ImmExt, PCTarget);
  mux2 #(32)  pcmux(PCPlus4, PCTarget, PCSrc, PCNext);

  // Register file and immediate generation
  regfile rf(clk, RegWrite, Instr[19:15], Instr[24:20], Instr[11:7], Result, SrcA, WriteData);
  extend ext(Instr[31:7], ImmSrc, ImmExt);

  // ALU logic
  mux2 #(32)  srcbmux(WriteData, ImmExt, ALUSrc, SrcB);
  alu         alu(SrcA, SrcB, ALUControl, ALUResult, Zero);
  mux3 #(32)  resultmux(ALUResult, ReadData, PCPlus4, ResultSrc, Result); 
  
  //// [MODIFICAÇAO] nessa linha onde agora tem PCPlus4, antes era 32'b0 (zero) o que nao tinha utilidade e fazia nao dar suporte a instruçoes de JAL
  //// agora é possivel fazer o jump e link, ou seja, guardar o endereco de retorno no registrador 
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module regfile(input  logic        clk, 
               input  logic        we3, 
               input  logic [ 4:0] a1, a2, a3, 
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0];

  // three ported register file
  // read two ports combinationally (A1/RD1, A2/RD2)
  // write third port on rising edge of clock (A3/WD3/WE3)
  // register 0 hardwired to 0

  always_ff @(posedge clk)
    if (we3) rf[a3] <= wd3;	

  assign rd1 = (a1 != 0) ? rf[a1] : 0;
  assign rd2 = (a2 != 0) ? rf[a2] : 0;
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


module adder(input  [31:0] a, b,
             output [31:0] y);

  assign y = a + b;
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module extend(input  logic [31:7] instr,
              input  logic [1:0]  immsrc,
              output logic [31:0] immext);

  assign immext = 
    (immsrc == 2'b00) ? {{20{instr[31]}}, instr[31:20]} : // I-type  //// [MODIFICAÇAO] formato I-Type adicionado
    //// Adicionado para dar suporte para instruçoes aritimeticas com imediato e instruçoes de load

    (immsrc == 2'b01) ? {{20{instr[31]}}, instr[31:25], instr[11:7]} : // S-type
    
    (immsrc == 2'b10) ? {{20{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0} : // B-type //// [MODIFICAÇAO] formato B-Type adicionado
    //// Bits reorganizados em B-Type para fazer corretamente o calculo do offset para o endereco do branch
                        //extensao sinal | bit 12 | bit 11 | bits 10-5 | bits 4-1 | bit 0
    
    (immsrc == 2'b11) ? {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0} : // J-type
    32'bx; // default
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module flopr #(parameter WIDTH = 8)
              (input  logic             clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module mux2 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, 
              input  logic             s, 
              output logic [WIDTH-1:0] y);

  assign y = s ? d1 : d0; 
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module mux3 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, d2,
              input  logic [1:0]       s, 
              output logic [WIDTH-1:0] y);

  assign y = s[1] ? d2 : (s[0] ? d1 : d0); 
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module imem(input  logic [31:0] a,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0];

  initial
      $readmemh("riscvtest.txt",RAM,0 , 20);

  assign rd = RAM[a[31:2]]; // word aligned
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module dmem(input  logic        clk, we,
            input  logic [31:0] a, wd,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0];

  assign rd = RAM[a[31:2]]; // word aligned

  always_ff @(posedge clk)
    if (we) RAM[a[31:2]] <= wd;
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module alu(input  logic [31:0] a, b,
           input  logic [2:0]  alucontrol,
           output logic [31:0] result,
           output logic        zero);

  logic [31:0] condinvb, sum;
  logic        v;              // overflow
  logic        isAddSub;       // true when is add or subtract operation

  assign condinvb = alucontrol[0] ? ~b : b;
  assign sum = a + condinvb + alucontrol[0];
  assign isAddSub = ~alucontrol[2] & ~alucontrol[1] |
                    ~alucontrol[1] & alucontrol[0];

  assign result = 
    (alucontrol == 3'b000) ? sum :              // add
    (alucontrol == 3'b001) ? sum :              // sub  
    (alucontrol == 3'b010) ? (a & b) :          // and
    (alucontrol == 3'b011) ? (a | b) :          // or  
    (alucontrol == 3'b100) ? (a ^ b) :          // xor
    (alucontrol == 3'b101) ? (sum[31] ^ v) :    // slt
    (alucontrol == 3'b110) ? (a << b[4:0]) :    // sll
    (alucontrol == 3'b111) ? (a >> b[4:0]) :    // srl
    32'bx;

  assign zero = (result == 32'b0);
  assign v = ~(alucontrol[0] ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;
  
endmodule